grammar edu:umn:cs:melt:exts:ableC:parallel:impl:bthrdpool;

marking terminal BThrdpool_t 'bthrdpool' lexer classes {Keyword, Reserved};

concrete productions top::TypeQualifier_c
| 'bthrdpool' {
    top.typeQualifiers = foldQualifier([bthrdpoolParallelQualifier(location=top.location)]);
    top.mutateTypeSpecifiers = [];
  }

abstract production bthrdpoolParallelQualifier
top::Qualifier ::=
{
  top.pp = text("bthrdpool");
  top.mangledName = "bthrdpool";
  top.qualIsPositive = true;
  top.qualIsNegative = false;
  top.qualAppliesWithinRef = true;
  top.qualCompat = \qtc::Qualifier ->
    case qtc of bthrdpoolParallelQualifier() -> true | _ -> false end;
  top.qualIsHost = false;
  top.errors := [];

  top.parSystem = just(bthrdpoolParallelSystem());
}
