grammar edu:umn:cs:melt:exts:ableC:parallel:concretesyntax;

marking terminal Spawn_t 'spawn' lexer classes {Keyword, Reserved};
marking terminal Sync_t 'sync' lexer classes {Keyword, Reserved};
marking terminal Parallel_t 'parallel' lexer classes {Keyword, Reserved};

terminal By_t 'by' lexer classes {Keyword, Reserved};
terminal As_t 'as' lexer classes {Keyword, Reserved};
terminal In_t 'in' lexer classes {Keyword, Reserved};
