grammar edu:umn:cs:melt:exts:ableC:parallel:exts:balancer;

exports edu:umn:cs:melt:exts:ableC:parallel:exts:balancer:base;
