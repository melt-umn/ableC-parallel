grammar edu:umn:cs:melt:exts:ableC:parallel;

exports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:parallel:concretesyntax;
