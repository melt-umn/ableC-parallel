grammar edu:umn:cs:melt:exts:ableC:parallel:impl:bworkstlr;

imports edu:umn:cs:melt:ableC:concretesyntax;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports edu:umn:cs:melt:ableC:abstractsyntax:overloadable;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:balancer;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:parallel;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:parallel:loop;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:parallel:spawn;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:sync;

imports edu:umn:cs:melt:exts:ableC:parallel:impl:workstlr;

imports edu:umn:cs:melt:exts:ableC:constructor:abstractsyntax;
