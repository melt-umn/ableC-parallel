grammar edu:umn:cs:melt:exts:ableC:parallel:exts:balancer:base;

imports edu:umn:cs:melt:ableC:concretesyntax;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;

imports edu:umn:cs:melt:exts:ableC:constructor:abstractsyntax;
