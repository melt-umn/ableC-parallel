grammar edu:umn:cs:melt:exts:ableC:parallel:exts:synchronization:abstractsyntax;

abstract production synchronizedType
top::ExtType ::= sys::LockSystem inner::Type sync::SynchronizationDesc
                  pp::Document mangledName::String
{
  propagate canonicalType;

  top.pp = pp;

  top.host = extType(top.givenQualifiers, refIdExtType(structSEU(), just(mangledName), 
    s"edu:umn:cs:melt:exts:ableC:parallel:exts:synchronization:${mangledName}"));
  top.mangledName = mangledName;
  top.isEqualTo =
    \ other::ExtType ->
      case other of
      | synchronizedType(_, _, _, _, mn) -> mn == mangledName
      | _ -> false
      end;

  -- Override new and delete to actually do important things
  top.newProd = 
    just(\e::Exprs l::Location -> synchronizedNew(e, top, location=l));
  top.deleteProd = just(\e::Expr -> synchronizedDelete(e, top));
  -- TODO: exprInitProd, objectInitProd (it would be nice to support these so
  -- we don't have to use the new ...(...), but the implementation is not
  -- incomplete without them

  -- Override literally everything else to make it an error
  local errExpr :: (Expr ::= Location) =
    \loc::Location -> errorExpr([err(loc, "A `synchronized` object cannot be accessed outside of a holding block")], location=loc);

  -- FIXME:
  -- Should some of these not be included? i.e. should we check whether
  -- these operations are even defined on the inner type?
  top.ovrld:arraySubscriptProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:callProd = just(\e::Expr es::Exprs l::Location -> errExpr(l));
  top.ovrld:callMemberProd = just(\e::Expr b::Boolean n::Name es::Exprs l::Location -> errExpr(l));
  top.ovrld:memberProd = just(\e::Expr b::Boolean n::Name l::Location -> errExpr(l));
  top.ovrld:preIncProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:preDecProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:postIncProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:postDecProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:addressOfArraySubscriptProd = just(\e::Expr i::Expr l::Location -> errExpr(l));
  top.ovrld:addressOfCallProd = just(\e::Expr h::Exprs l::Location -> errExpr(l));
  top.ovrld:addressOfMemberProd = just(\e::Expr b::Boolean n::Name l::Location -> errExpr(l));
  top.ovrld:dereferenceProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:positiveProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:negativeProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:bitNegateProd = just(\e::Expr l::Location -> errExpr(l));
  top.ovrld:notProd = just(\e::Expr l::Location -> errExpr(l));
  
  -- We have to allow this so we can allow constructions using 'new'
  top.ovrld:lEqProd = just(\x::Expr r::Expr l::Location -> synchronizedLEq(x, r, 
                                  sys, sync, mangledName, location=l));
  
  top.ovrld:rEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:eqArraySubscriptProd = just(\e::Expr i::Expr x::Expr l::Location -> errExpr(l));
  top.ovrld:eqCallProd = just(\e::Expr a::Exprs x::Expr l::Location -> errExpr(l));
  top.ovrld:eqMemberProd = just(\e::Expr b::Boolean n::Name x::Expr l::Location -> errExpr(l));
  
  top.ovrld:lMulEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rMulEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lDivEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rDivEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lModEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rModEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lAddEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rAddEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lSubEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rSubEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lLshEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rLshEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lRshEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rRshEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lAndEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rAndEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lXorEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rXorEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lOrEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rOrEqProd = just(\x::Expr r::Expr l::Location -> errExpr(l));

  top.ovrld:lAndProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rAndProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lOrProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rOrProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  
  top.ovrld:lAndBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rAndBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lOrBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rOrBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  
  top.ovrld:lXorProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rXorProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  
  top.ovrld:lLshBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rLshBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lRshBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rRshBitProd = just(\x::Expr r::Expr l::Location -> errExpr(l));

  top.ovrld:lEqualsProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rEqualsProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lNotEqualsProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rNotEqualsProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  
  top.ovrld:lLtProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rLtProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lGtProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rGtProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lLteProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rLteProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lGteProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rGteProd = just(\x::Expr r::Expr l::Location -> errExpr(l));

  top.ovrld:lAddProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rAddProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lSubProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rSubProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lMulProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rMulProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lDivProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rDivProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:lModProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
  top.ovrld:rModProd = just(\x::Expr r::Expr l::Location -> errExpr(l));
}
  
abstract production synchronizedLEq
top::Expr ::= l::Expr r::Expr sys::LockSystem desc::SynchronizationDesc
              mangledName::String
{
  top.pp = ppConcat([l.pp, space(), text("="), space(), r.pp]);
  forwards to 
    case r of
    | newExpr(_, consExpr(arg, nilExpr())) ->
        initializeSynchronized(l, arg, sys, desc, mangledName, location=top.location)
    | newExpr(_, _) -> errorExpr(
        [err(top.location, "A `synchronized` object should be constructed from a single argument")],
        location=top.location)
    | _ -> errorExpr(
      [err(top.location, 
        "A `synchronized` object cannot be accessed outside of a holding block")],
      location=top.location)
    end;
}

abstract production synchronizedNew
top::Expr ::= e::Exprs syncType::ExtType
{
  top.pp = ppConcat([text("new"), space(), syncType.pp, 
    parens(ppImplode(comma(), e.pps))]);

  forwards to
    errorExpr([err(top.location,
      "Construction of a `synchronized` object only allowed on the rhs of an assignment")],
      location=top.location);
}

abstract production initializeSynchronized
top::Expr ::= l::Expr ex::Expr sys::LockSystem desc::SynchronizationDesc
              mangledName::String
{
  top.pp = ppConcat([lhs.pp, text(" = "), ex.pp]);

  local lhs::Expr = exprAsType(l,
    extType(nilQualifier(),
      refIdExtType(structSEU(), just(mangledName),
        s"edu:umn:cs:melt:exts:ableC:parallel:exts:synchronization:${mangledName}")),
    location=top.location);

  lhs.env = top.env;
  lhs.controlStmtContext = top.controlStmtContext;

  forwards to
    ableC_Expr {
      ({
        $Expr{lhs}.value = $Expr{ex};
        $Expr{sys.initializeLock(ableC_Expr{$Expr{lhs}.lck}, nilExpr(), top.location)};

        $Stmt{foldStmt(map(
          \p::Pair<String Pair<Boolean Expr>> ->
            ableC_Stmt { 
              $Expr{sys.initializeCondvar(
                ableC_Expr{$Expr{lhs}.$name{if !p.snd.fst then s"__not__${p.fst}" else s"__${p.fst}"}},
                  consExpr(
                    explicitCastExpr(
                      typeName(
                        extTypeExpr(nilQualifier(), lockType(sys)),
                        pointerTypeExpr(nilQualifier(),
                          baseTypeExpr())
                      ),
                      ableC_Expr{&($Expr{lhs}.lck)},
                      location=top.location
                    ),
                    nilExpr()
                  ),
                  top.location
                )};
            },
          desc.conditions))}
        
        $Expr{lhs};
      })
    };
}

abstract production synchronizedDelete
top::Stmt ::= e::Expr syncType::ExtType
{
  top.pp = ppConcat([text("delete"), space(), e.pp]);

  local sys::LockSystem =
    case syncType of
    | synchronizedType(s, _, _, _, _) -> s
    | _ -> error("This function only called by being this type")
    end;
  local desc::SynchronizationDesc =
    case syncType of
    | synchronizedType(_, _, d, _, _) -> d
    | _ -> error("This function only called by being this type")
    end;

  sys.env = top.env;

  forwards to
    ableC_Stmt {
      {
        struct $name{syncType.mangledName}* __obj = 
          (struct $name{syncType.mangledName}*) &$Expr{e};
        $Stmt{sys.lockDeleteProd.fromJust(ableC_Expr{&(__obj->lck)})}
        $Stmt{foldStmt(map(
          \p::Pair<String Pair<Boolean Expr>> ->
              sys.condvarDeleteProd.fromJust(
                ableC_Expr{&(__obj->$name{if !p.snd.fst then s"__not__${p.fst}" else s"__${p.fst}"})}
              ),
          desc.conditions
        ))}
      }
    };
}
