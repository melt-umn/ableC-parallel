grammar edu:umn:cs:melt:exts:ableC:parallel:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports silver:langutil only ast;

imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;

