grammar edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;

global builtin :: Location = builtinLoc("parallel");
