grammar well_definedness;

{-  This silver specification does not generate a useful working
    compiler, it only serves as a grammar for running the modular
    well-definedness analysis. -}

import edu:umn:cs:melt:ableC:host;
import edu:umn:cs:melt:exts:ableC:parallel:impl:vector;
