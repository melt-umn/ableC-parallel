grammar edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:spawn;

imports edu:umn:cs:melt:ableC:abstractsyntax:host;
