grammar edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:parallel;

imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:parallel:loop;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports edu:umn:cs:melt:exts:ableC:constructor:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp;
