grammar edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax:locks;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:exts:ableC:constructor:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;
