grammar edu:umn:cs:melt:exts:ableC:parallel:exts:synchronization:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports edu:umn:cs:melt:exts:ableC:parallel:exts:synchronization:abstractsyntax;

imports silver:langutil;
