grammar edu:umn:cs:melt:exts:ableC:parallel:exts:balancer:impl:fcfs;

imports edu:umn:cs:melt:ableC:concretesyntax;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports edu:umn:cs:melt:ableC:abstractsyntax:overloadable as ovrld;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:exts:ableC:parallel:abstractsyntax;
imports edu:umn:cs:melt:exts:ableC:parallel:exts:balancer;

imports edu:umn:cs:melt:exts:ableC:constructor:abstractsyntax;
