grammar determinism;

import edu:umn:cs:melt:ableC:host only ablecParser;

copper_mda testConcreteSyntax(ablecParser) {
  edu:umn:cs:melt:exts:ableC:parallel:concretesyntax;
}

